*
* diodes.lib
*

* Some diode models to test if reading Spice libraries works.

* Not really 1N4148, just shoddily based on some values in datasheet.
.MODEL 1N4148 D (BV=100 CJO=4p IBV=100u IS=4n M=0.33 N=2
+ RS=0.5 TT=10n VJ=0.8)

* The below models have made up values - I didn't bother to check if they are physically correct.


.model D1 D(Is=1.23n N=1.23 Rs=.7890 Ikf=12.34m Xti=3 Eg=1.23 Cjo=.90p
+           M=.56 Vj=.78 Fc=.9 Isr=12.34n Nr=2.345 Bv=100 Ibv=100u Tt=12.34n)

* This line has a single trailing space.
* DUsual* models always have the same values to save space on test asserts.
.model D2_Usual D(BV=1.1U CJO=2.2M IBV=3.3 IS=4.4K M=5.5MEG N=6.6G) 

* Trailing spaces, and an (empty) continuation.
.model D3_Usual D(BV=1.1U CJO=2.2M IBV=3.3 IS=4.4K M=5.5MEG N=6.6G 
+) 

.model D4  D( Is=0.1p 
+             Rs=2 
+             CJO=3p 
+             Tt=45n ; Test comment
+             Bv=678 
+             Ibv=0.1p )
* (Has trailing spaces after each parameter value)

.model D5_Empty D () ; Empty model

* Parentheses are optional.
.model D6_Empty D

.model D7_Empty D ; Empty model, no parentheses, ending with a comment.

.model D8_Empty D

.model D9_Empty D;

* Several parameters, no parentheses.
.model D10_Usual D BV=1.1U CJO=2.2M IBV=3.3 IS=4.4K M=5.5MEG N=6.6G

* Several parameters, no parentheses, multiple lines.
.model D11_Usual D BV=1.1U
+                  CJO=2.2M
+                  IBV=3.3;
+                  IS=4.4K ; Test comment
+                  M=5.5MEG
+                  N=6.6G

.model D12_Usual D
+BV=1.1U 
+CJO=2.2M 
+IBV=3.3;
+IS=4.4K;
+M=5.5MEG 
+N=6.6G 

* Test some parameter synonyms.
.model D13_Usual D
+ BV=1.1U
+ CJ0=2.2M
+ IBV=3.3
+ JS=4.4K
+ MJ=5.5MEG
+ N=6.6G
.model D14_Usual D
+ BV=1.1U
+ CJ=2.2M
+ IBV=3.3
+ JS=4.4K
+ MJ=5.5MEG
+ N=6.6G

* Two spaces as a separator everywhere, two trailing spaces.
.model  D15_Usual  D  (  BV=1.1U  CJ=2.2M  IBV=3.3  JS=4.4K  MJ=5.5MEG  N=6.6G  )  

* Spaces aligning param names and values.
.model D16_Usual D
+ BV  = 1.1U
+ CJ0 = 2.2M
+ IBV = 3.3
+ JS  = 4.4K
+ MJ  = 5.5MEG
+ N   = 6.6G

* No newline at the end of file.
.model D17_Usual D(BV=1.1U CJ=2.2M IBV=3.3 JS=4.4K MJ=5.5MEG N=6.6G)
