.title KiCad schematic
.include "diodes.lib"
.tran 1u 10m

C1 /out GND 10u
R1 /out GND 100k
D1 /in /out DIODE1
V1 /in GND SIN( 0 5 10k    )
.end
